module Out_s2(

);
endmodule