`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 08.07.2025 06:20:59
// Design Name: 
// Module Name: NeuronROM
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module NeuronROM(
    output logic signed [34:0] Weights1 [143:0],
    output logic signed [34:0] Weights2 [143:0],
    output logic signed [34:0] Weights3 [143:0],
    output logic signed [34:0] Weights4 [143:0]
    );

    always_comb begin
        Weights1= '{35'sh1CA2E6C00, 35'shFC95B6CC0, 35'shF01D4E000, 35'shC3539100 , 35'shAC43350  , 35'shE7F29E600, 35'shF414EAC00, 35'shE8F27F00, 35'shE39AF7C00, 35'shED6211400, 35'shFB61BD300, 35'shFB2297100, 35'shDE3D08400, 35'sh79E6A480, 35'shF94C44E80, 35'sh12C6F0E00, 35'shD4074B000, 35'shF6E3AA700, 35'sh851D4A00, 35'sh1778D6A00, 35'shE6F74CC00, 35'shF89030100, 35'shB773ED00, 35'sh506DE600, 35'shF3464F400, 35'shE4E845000, 35'shA6939600, 35'sh8E7B3B00, 35'shE1E678A00, 35'shFF9282588, 35'shE07AEFC00, 35'shF80F29F00, 35'shD031FC000, 35'shF53B3E500, 35'shAE3709, 35'shB2E94F00, 35'shEB5494E00, 35'shF13184500, 35'sh9FA27700, 35'sh6EFBCE00, 35'shD08168C00, 35'sh60CCB800, 35'sh802D3300, 35'sh187274400, 35'shD3F710800, 35'shC0941800, 35'shF20F30500, 35'sh3D87854, 35'shF48CE6700, 35'shFBDC35700, 35'shDA74FC400, 35'shFBC00C700, 35'sh1ADDF1A0, 35'shFB754D880, 35'shEFA731200, 35'shEA804600, 35'shE31E12000, 35'shF4D3DB400, 35'shE1C83B400, 35'sh89C69600, 35'shE3A046A00, 35'sh9B763900, 35'shFB38DDD80, 35'sh106781000, 35'shE23AC2800, 35'shED0B49E00, 35'sh457D9500, 35'sh4DBD2C00, 35'shF620A9B00, 35'shA06EE100, 35'shE49CED600, 35'sh256D65400, 35'shD66EA3000, 35'shB8CF3500, 35'shFEF688C60, 35'shFE0F95880, 35'shFAF488B00, 35'sh10EBF1400, 35'shEF32F1600, 35'shF5816D00, 35'shE0D588A00, 35'shF89AA8D00, 35'shF927D6480, 35'sh197787200, 35'shE8008E200, 35'shEAE620400, 35'shEC5A3500, 35'shFE40EAE40, 35'shF821C5E80, 35'sh12E50F000, 35'shFDFFD200, 35'sh74B9ED00, 35'shDB7213C00, 35'sh83555200, 35'shEF7CDD200, 35'sh7B808080, 35'shDFF4BBC00, 35'shBDDA5900, 35'shEDB64EA00, 35'sh9C8A2900, 35'shD7D259400, 35'sh52CDB800, 35'shE1003F400, 35'sh1B1C4D200, 35'shE127AAA00, 35'sh11F26BA00, 35'sh10C93A400, 35'sh16324EC00, 35'sh950FDB00, 35'shFAB568180, 35'shE9C10AA00, 35'sh22F8A2400, 35'shFC9B81E00, 35'sh53CB4480, 35'shF9F45CA80, 35'sh10CF50E00, 35'shEEFD88C00, 35'shFE7E62640, 35'shF6C80AE00, 35'sh1AF8DD800, 35'shFBF5E0F80, 35'sh77325180, 35'shFCDCDE900, 35'sh117D9CE00, 35'shF7EF85400, 35'sh104EF9600, 35'shE5AA1E400, 35'sh2152A640, 35'shB10D9200, 35'sh1133CE400, 35'shFDBD1B440, 35'sh18F8E7400, 35'shF67B66400, 35'shF4017EF00, 35'shF1F67AD00, 35'sh7C60F58, 35'shF16781100, 35'sh28A6938, 35'shF9696B800, 35'shEA7DE800, 35'shEE7412000, 35'sh196945800, 35'shE688ECE00, 35'shFD0B21B00};
        Weights2= '{35'shC1D808000, 35'shFF9CC9DA0, 35'shDE0779C00, 35'sh17B34B600, 35'shDA7A1DC00, 35'shF44DE1E00, 35'sh1A083F200, 35'sh1473D8400, 35'sh22296780, 35'shF16043D00, 35'shF341CB100, 35'shFEEA7F220, 35'sh19C15C600, 35'shFEB8AD840, 35'shF0AF2D200, 35'sh50C81B80, 35'shB5A51300, 35'shEEDA51400, 35'shEEB74C200, 35'sh76FBC10, 35'shEBA53100, 35'shF5D2AC800, 35'shF61B74F00, 35'shF4A4C3B00, 35'shCDFD9EC00, 35'sh10343CA00, 35'shF7CCC7F00, 35'sh152A0C000, 35'shECFD12400, 35'shFC82A600, 35'sh60A87F80, 35'shFE68DFB20, 35'shF9C6AF000, 35'shF49C24800, 35'sh33553F80, 35'sh51D03D80, 35'shF859B5A00, 35'sh106355C00, 35'sh1C050000, 35'sh11AC71A00, 35'shEB0C55200, 35'shFE7895440, 35'sh86420200, 35'shEABC4100, 35'shE8A54D600, 35'sh10E4C660, 35'sh57B31380, 35'sh35B9DDC0, 35'shDD3F04400, 35'sh2B8A83400, 35'shF429C0600, 35'sh200C6E400, 35'sh5EEA4780, 35'sh51B06980, 35'shE0F18B00, 35'sh14983B600, 35'shF823CD00, 35'sh10A96A800, 35'sh285E8E000, 35'sh921FA700, 35'sh114598E00, 35'sh2141D9000, 35'sh100E83800, 35'shF5F34EE00, 35'shF89584680, 35'sh275CDC40, 35'sh9710A300, 35'sh21843B40, 35'shFA35E0B00, 35'sh15186A000, 35'shF6FC23F00, 35'sh13FA82200, 35'shAB0E8200, 35'sh27352A800, 35'sh11D465000, 35'sh193979E0, 35'shF603E1D00, 35'sh1F85CDE00, 35'sh146E9C400, 35'shA9EDBF00, 35'sh84CF6100, 35'shFF3F392F0, 35'sh119E9EE00, 35'sh57329800, 35'sh1DCE72E00, 35'sh60C9D680, 35'sh22F671800, 35'sh277D08C0, 35'shFFFD9850C, 35'sh178B1F600, 35'sh626D5780, 35'shFC563B5C0, 35'shD680DB00, 35'sh173488600, 35'shF5BF5CF00, 35'shF70E48A00, 35'shF2D647800, 35'shE9054700, 35'shF6DAABC00, 35'shF84948F00, 35'shF800D3C80, 35'shFF097DB30, 35'sh1CC51D000, 35'sh57FCD900, 35'sh240972C00, 35'shFD577A400, 35'sh108F0AA00, 35'sh47E4E380, 35'shFB1EA8A80, 35'sh19AE4E800, 35'sh1666CC400, 35'sh117EC2800, 35'sh33C96400, 35'shFC0401C40, 35'sh12941FE00, 35'shEFFA1E400, 35'sh4CA21100, 35'shFFDB6EC84, 35'sh1F944A400, 35'sh10A8B9400, 35'sh12F7CB800, 35'sh10EE52000, 35'sh150520800, 35'shFBE611A00, 35'sh16BE5DC00, 35'sh169658200, 35'shEF8CBD00, 35'shF96740B80, 35'shFFDC6641C, 35'shF3A86FB00, 35'shFC3453580, 35'sh10DC23500, 35'sh18B4D9200, 35'shF12BFC900, 35'shF4EC6E200, 35'sh59174680, 35'shCB87EC00, 35'shFDD48DC00, 35'sh195BA7C00, 35'sh9BE4E700, 35'shF826D3D00, 35'sh42D63F00, 35'sh1AC9B0000, 35'shE9FE23000};
        Weights3= '{35'sh8EA2F100 , 35'shF23C5DF00, 35'sh1C7AC3C00, 35'shD86BCA400, 35'sh1AF48FC00, 35'shECE65EC00, 35'shCABAD500, 35'shFB673CC80, 35'shFB2977E80, 35'shF9059AA80, 35'sh130915A00, 35'shFD6CA5040, 35'sh20B839C00, 35'shF99902980, 35'sh1BDE79200, 35'sh5CDED800, 35'sh1FD729400, 35'shE3FF48800, 35'sh4644098, 35'shF15FF2F00, 35'sh12F0A9E00, 35'shD9E786800, 35'sh15A3C2E00, 35'shF161CF100, 35'sh61830E00, 35'shEF6EBA000, 35'sh19EEBB800, 35'shE6AB70A00, 35'sh134B79600, 35'shE637B6A00, 35'sh4F505880, 35'shDB5EA4000, 35'shFFE066E68, 35'sh10519AE00, 35'shD78D3C00, 35'shF90275200, 35'sh115BF7E00, 35'sh13AD82C00, 35'shB25EDF00, 35'shF84168D00, 35'shF0A5BC00, 35'shED7F79C00, 35'sh15088EE00, 35'shDC2177C00, 35'sh295D6500, 35'shF09635200, 35'shF20E0AC00, 35'shDE87C5C00, 35'shF094FFB00, 35'shF74875600, 35'shEE5B2200, 35'shE05CA0600, 35'shF513C3700, 35'shEC0AD5200, 35'shEC4D1600, 35'shE2E7FF600, 35'sh10780E200, 35'shED3034200, 35'sh13957D800, 35'shE3A3DA200, 35'shF4BBCBC00, 35'shC686FA00, 35'shFA3E5FF80, 35'shFC731DDC0, 35'sh191908200, 35'sh4DCB0600, 35'sh1183D1000, 35'shD81B2BC00, 35'shEEFF4F600, 35'shE64883C00, 35'shEF933C600, 35'shD89548C00, 35'shFAD9FEF00, 35'shDD9CB3000, 35'shFA0CB9B80, 35'shF5791DE00, 35'sh4C22F700, 35'shFA814A400, 35'shF40B87000, 35'shDE12FC800, 35'shF8FD55700, 35'shF86693500, 35'sh193593500, 35'sh6E81DA80, 35'sh22610F40, 35'shFB7701D00, 35'sh18DC2BE00, 35'shFA58BD880, 35'shF7BAE2C00, 35'shE33AEF200, 35'sh9B8A5C00, 35'shE657BF400, 35'shDC2F3100, 35'shE885D8A00, 35'sh13FBE2400, 35'shFE877BDC0, 35'sh9D166800, 35'shE6B09F400, 35'sh174F8EE00, 35'shB339210, 35'sh200082800, 35'shE2596FE00, 35'sh4001B600, 35'shE7BD2CE00, 35'sh26B77AC00, 35'shEC9243E00, 35'shF90D48800, 35'shF5A37A700, 35'shB1A46A00, 35'shE1380FC00, 35'sh1A5DF2400, 35'shDB5234800, 35'sh1A1DB1C00, 35'shF9DF72880, 35'sh13FCD5600, 35'shDDDF44C00, 35'shFC12F64C0, 35'sh19C03760, 35'shFDD82DA00, 35'shFF92B8848, 35'sh2582F6400, 35'shFAF30D180, 35'sh140D35000, 35'shE47E88000, 35'sh1FE9DD800, 35'shE34BB9E00, 35'sh21BF70400, 35'shDAE14C400, 35'sh295C1D40, 35'shE3E95BA00, 35'sh18766C400, 35'shD257C4800, 35'sh1BDDCC600, 35'shDE4F11400, 35'shFD9234900, 35'shF8244F380, 35'shD4DC3A00, 35'shFAE4BE380, 35'shC37FE400, 35'shF0C011800, 35'sh9BD2F20, 35'sh3CC49140, 35'sh1EB89C200, 35'shDD1E71C00};
        Weights4= '{35'sh273B64C00, 35'sh2E7AB8800, 35'sh9708D000 , 35'shEC018B400, 35'sh1E4284A00, 35'shA1678300, 35'shF1BC3A500, 35'shEC6E7EE00, 35'sh16E54FC00, 35'shFAC21E00, 35'shF5703D200, 35'shFBCE08C00, 35'sh17B08A400, 35'sh93766700, 35'shF7DA8A800, 35'shF805A5180, 35'shF41387300, 35'sh1EC80A600, 35'shD1882300, 35'shFDD86E00, 35'shF5D610D00, 35'sh2024E2800, 35'sh967B5D00, 35'shF7E3ED000, 35'sh1C07C8200, 35'sh439ED580, 35'sh209C8D40, 35'shFE1D71560, 35'sh16227D800, 35'sh11AAA2A00, 35'sh50009080, 35'sh3C3267C0, 35'shFE8072080, 35'shC6D3980, 35'shF75740A00, 35'shB3DA4500, 35'sh1ECD58800, 35'shEF214F800, 35'shEE63BFE00, 35'sh1A35B6A00, 35'sh1DC759000, 35'sh84E92700, 35'shF68340A00, 35'shFED192FC0, 35'sh26A499000, 35'sh18CB21200, 35'sh58E89380, 35'shFAC44800, 35'sh115581200, 35'shE59781400, 35'shE8DBA100, 35'shE1E1EFE00, 35'sh1318E6400, 35'shE45146600, 35'shF9D0C9300, 35'shF624A1300, 35'shF3BEC2300, 35'shCE901100, 35'shE77D6BC00, 35'shF45721300, 35'shE80A23200, 35'sh46224E00, 35'sh58602B00, 35'sh2A03FA00, 35'shFDE19C100, 35'shF990D8680, 35'shF98810000, 35'shE44850A00, 35'sh25B73B80, 35'sh6834BA80, 35'sh4A1EB980, 35'sh6663C500, 35'sh271BB5400, 35'shD1D6B5C00, 35'sh4C406100, 35'shFCE66B1C0, 35'shC6C9A300, 35'sh158BAD60, 35'shF5AC4800, 35'shAD89FC0, 35'shE332C1400, 35'shF9B9A0180, 35'shE443DB600, 35'shF59F33300, 35'shF5F9EDB00, 35'shF9C835F80, 35'shEA07A2E00, 35'shEF32ABA00, 35'sh29A84180, 35'shFEF753520, 35'shA71A4000, 35'shEACEF4400, 35'shE72E19600, 35'shE26FD2E00, 35'shFC408A540, 35'shFE1A90800, 35'shF4BAF4A00, 35'shE5281FA00, 35'sh9F70C700, 35'sh178E8480, 35'shF43AAFA00, 35'shF518FFD00, 35'shE44AD6400, 35'shFE3249160, 35'shFF78B4510, 35'sh181035E00, 35'shF72895B00, 35'sh6A47690, 35'shD6FA1F800, 35'shF2D6D0900, 35'shE86918200, 35'sh1C5000000, 35'shF10038400, 35'sh448A2B00, 35'sh518F7180, 35'sh125DC9400, 35'shEBE4EB800, 35'shE0EEB4600, 35'shF49642300, 35'sh98BDC000, 35'shF09E78E00, 35'shF25C7DC00, 35'sh7E873B80, 35'sh12B469A00, 35'shFD537B880, 35'sh1CA1E3800, 35'sh81516700, 35'sh77929F00, 35'shDF172C800, 35'shFA2CD4980, 35'shD51F73000, 35'shA271F400, 35'shE7757E600, 35'sh2F358840, 35'shE5FBF8200, 35'sh83C51900, 35'shD40AF5800, 35'shEF0875C00, 35'shE7163A600, 35'shFBD0DC380, 35'shE3738E000, 35'sh1035EEC00, 35'sh219271C0, 35'sh3FAF0F00};
    end

endmodule
