


module Filtros_s2_ROM#
(
    parameter WIDTH = 17
)
(
    //FiltroX = [Fila][Columna][Canal] (es más simple la multiplexación escrita de esta manera)
    //input logic[WIDTH-1:0]  F1[2:0][2:0][2:0],
    //input logic[WIDTH-1:0]  F2[2:0][2:0][2:0],
    //input logic[WIDTH-1:0]  F3[2:0][2:0][2:0],

    output logic signed [WIDTH-1:0] Filtro1[2:0][2:0][2:0],
    output logic signed [WIDTH-1:0] Filtro2[2:0][2:0][2:0],
    output logic signed [WIDTH-1:0] Filtro3[2:0][2:0][2:0],
    output logic signed [WIDTH-1:0] Filtro4[2:0][2:0][2:0]
);
    always_comb begin
        // Filtro1[canal][COLUMNA][fila] - Formato Q0.16 (1 bit de signo, 16 bits fraccionales)
    Filtro1 = '{
  '{ // Canal 0
    '{17'sb1110101101011110, 17'sb1101010111010000, 17'sb1011010100101001}, // Columna 0: Filas 0,1,2
    '{17'sb1101100110111101, 17'sb1110010010000101, 17'sb1101101011000000},
    '{17'sb1111001000110110, 17'sb1111100011101001, 17'sb1110010001111101}
  },
  '{ // Canal 1
    '{17'sb1110100001011111, 17'sb0000111001101101, 17'sb0101010011101001},
    '{17'sb1110110001101110, 17'sb1111010000100101, 17'sb0100010100000000},
    '{17'sb1111001000010011, 17'sb1111111110111000, 17'sb0100000000101110}
  },
  '{ // Canal 2
    '{17'sb1111110101101110, 17'sb1111100011000001, 17'sb1111101001100111},
    '{17'sb1111100111000001, 17'sb0011110111110101, 17'sb1111101100100101},
    '{17'sb1111110101101100, 17'sb1110101111111011, 17'sb0000011010000111}
  }
};

    Filtro2 = '{
  '{ // Fila 0
    '{17'sb0100101001110101, 17'sb1110010100000111, 17'sb1111110111011000},
    '{17'sb0011001000011100, 17'sb1111011110111110, 17'sb0001001100011000},
    '{17'sb0011111101101100, 17'sb1110101100111010, 17'sb0010010000011101}
  },
  '{ // Fila 1
    '{17'sb0100110101110001, 17'sb0000010101011010, 17'sb0011101110111011},
    '{17'sb0011011000110101, 17'sb1111101100100110, 17'sb0011111110011000},
    '{17'sb0001111011000011, 17'sb1111001100110001, 17'sb0011000011010101}
  },
  '{ // Fila 2
    '{17'sb0011000111111010, 17'sb0000011101111001, 17'sb1111011011000010},
    '{17'sb0010011101110001, 17'sb0000111001111001, 17'sb0100010111110100},
    '{17'sb0000000000000111, 17'sb1111110011000001, 17'sb1111111111101100}
  }
};
    Filtro3 = '{
  '{ // Canal 0
    '{17'sb0000101100001110, 17'sb0010010011111111, 17'sb0011001110101011}, // Columna 0: Filas 0,1,2
    '{17'sb0011001000100010, 17'sb0011011101111001, 17'sb0010100011011000},
    '{17'sb0000010110100010, 17'sb1111000100111111, 17'sb1111000010000111}
  },
  '{ // Canal 1
    '{17'sb1111000011100100, 17'sb1110101010010111, 17'sb1110101010000100},
    '{17'sb0010110110111001, 17'sb1111111001011111, 17'sb1111100111110110},
    '{17'sb0000010101100111, 17'sb0011001110110010, 17'sb0001110100011110}
  },
  '{ // Canal 2
    '{17'sb1111000010000010, 17'sb1111000011010001, 17'sb1110111100111010},
    '{17'sb0000010111010000, 17'sb0010101001000100, 17'sb1111010001100101},
    '{17'sb1111101000010111, 17'sb0001000111111101, 17'sb1111000010111001}
  }
};

    Filtro4 = '{
  '{ // Canal 0
    '{17'sb0000101100010011, 17'sb1110111101011010, 17'sb0001100011010100}, // Columna 0: Filas 0,1,2
    '{17'sb1111101110101000, 17'sb1111001011111100, 17'sb1111101100100011},
    '{17'sb1111000010000001, 17'sb1111101000010111, 17'sb1111010010010110}
  },
  '{ // Canal 1
    '{17'sb0100010100011110, 17'sb0011101101010101, 17'sb0010111001111110},
    '{17'sb0100000010001011, 17'sb0011100100011001, 17'sb0010110000000010},
    '{17'sb0010110111001001, 17'sb0010111101110111, 17'sb0011010100010101}
  },
  '{ // Canal 2
    '{17'sb1111110000111110, 17'sb0000111011111001, 17'sb1111011010101111},
    '{17'sb1111101000111100, 17'sb0010011111111011, 17'sb0000110011111010},
    '{17'sb0100010001111100, 17'sb0001110010000111, 17'sb0010100101110111}
  }
};

    end

endmodule