module Top(
    
);


endmodule